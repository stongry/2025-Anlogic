`protect begin_protected
`protect version = 1
`protect encrypt_agent = "Anlogic"
`protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-002"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
fwDAfTNMN7zICdZ5GlBN0t3S6ufLmVxeOb3CAp6eIqTNnUjCaJ4QJlT9Mrus24xB
a7KsbT2SmT/12lXpZwhxKnNqchTmewTW2vfKnHuhW+nt1g6/crLXR3RmSnsRlJWL
rUz778HdPZeVxxgwdSaCsgNhOy3OoKeW9DcmDOYoBXw=
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`protect key_block
fj84zIBrR1qdZpr/8sp8ja0ez8x7UJ7gqD9q+DO+nu0Pl8z9l1jaxX+J9TQ0L9iX
lieDNsvNm3bbMK5WVZxZfakrZ+OmGHzl5Yr6HZfqCgif/7eF/iN4KD09/AhweCRw
qohirS4dDVHrs9aFG7lRqcWqBMLYDpj6HFEncrLG/U4Y6yd9R63SrGq3NnCtJ/iv
Wrq9B3JOzuOs2aEriXLxvFLlZTTKXG7B9KILeqW1BX1/Rh1ThJ4j9IH0PAxIciQR
tH/WEQCopZC06BGO9pbuyxCwFov3D76BNvMEUU+DLhn74j5GPPeKvP4tkLQFO7Dq
S1hswlPNHJB9Y+uPQGETLA==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
fV9xjugOb0ROei46ce4Jr89zxlgtZjW9emWnEr63BT+SvrZfk7XA9IgV2EgapT0j
J0Kdiyfu8IWgmIjxCWeI7l9yotDIOLab6rAZtJ7GcRIO4LzvwAeThLo3CZCtoUrc
OoW66UX6HDFeK3MC6bqIG0u4Lo8fFt/Mo7lHxXC05RQ=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`protect key_block
e01A0xmn2UrGTKpahEEUwr3C8w1bP7MEY4xGJarn/ufqldH6XJVSb4oOJ8IA7Fmx
HJau8z3Bqq5olSryRo03fXh+TbOfEJoo0XChJ9I81AstVshYHGbW1KZ5LceFYodB
MtAfx6FxvDAIWUCgrX4+UUJYs5+piPbfj9IerYfjac16G8m2KYUENmJi9Rx9309r
/arC2oxx64Nd3zYThTwj2uJXcVZtjPtDv8CrXBxrmJtbSM6QUCSzMxHpoMDNILzP
gQIzFcEfTr40FdidoUyHSTw0jAmfW9CyWjoWCfUY0RwjR3eHKlX3ZjfAjglgw7+n
bMPoOdzfQgtWzH0PPnigeg==
`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
fYe5xNHJ/JNsJz2lr1QpA92t/VX8RrfXPyhsQaMCrhCyEb+6miNnXUuD/391b0fw
aQZkh5tm92nhUqVS2KsXzZxb8iuLaWAt134cSpnWQ/Z0tn9fi+LOdoW1sXOKA5zW
xAXBtZtQXhekd9tfTqgjrhi8zPiFo/FB/a3lMD0ATqs=
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 4128)
`protect data_block
TmJmOVhVYVpnU3c3eUZZYwDhH1Fcvg//nJ8V49hN6W/eWuwp5slRQ5ib/qKhrTAX
20mjIjZjeCypq2X7mnRMEaJbg2+4B/NWuNHTdm2WFRTyfUFAlRFaz9QT1TsBTU1+
1ZuEWbfUgl7Z6hq7Ww3aOhoDKlYuvjJ1GrNenIXUHZDmJ76clYYJiCUbQ1i2OKQb
uX9w+hBzjjsgKL4pxOVo2YcILleA9CkdYvOIxcJgrsYjEF+RAG3VHmXOKoUswX+J
+MDgv9l1J7hvd4VJPJvnETCsvgV0ImgFTgF73LwGH2qzmVQOdwJ/NZHU8hRhcXkp
2RsMdhrRkX7oPabkaqB7VSTOCTqzy/utFTrrGM8ije4nW2qsEIDBw5kwq0St3H8N
5rR+Zagq16Ttwy9YVJPwD8OKgEypdBmkcVuW/j09xHvmo7Jb6OdZxilfGoLHI1Ke
FfYvEcB5wn0MpvMbkGtVPcsAAkJaMiDL780kkF1aR7bOWmU5ajjE5ixXiRVljdT/
XqbQNY9CNxWdp1gJSbjtUBKdSJf01EoBHasti9N5EXfbkmyz3aIUvXVeprTsYEq4
NC0ux7ARJxILtWwOIjCRGK47rvB6Ow6ehJx3jK5mLJuarAtMagIxfE+WB8uEpjK/
j8s20G46kQhd2k1wVi6+ivEX52cRK4lA7z4uFOceMSr5abkqXpKBjgV8afdeSdso
QDmTdreltBVxYwUmB+Lf6eunWq98hxEpSN+wPlSMtA9iNyq3A7sL/d3Kh6a9Bm04
Jz6LhdGhubd3lCq4fQz/Zbj203BtQzsxVyXvHQ2V7tGVitxDsU1o+9Cvwp7SigIL
UJxhMcU1m1968M7Xq492GyS+qSDpwx8JtR7elx1KF0HdXoRiUPLdvWVRyvepYhr7
8ggyUdgUh41JVwvJJVwzwVtcaRygx8I5Klkte7MvQXvvc91B+HXum63aoCWj0OGd
da/NAZt45oTwbr35Q/E7xoFN+n+d0L4xHxp08pjPi7Jue9kUdL5GE54iK7T6K4Ph
UxgmqUuR1J5Z/8D6pj3La4rnR8sLWWXr+J7quDsTUY5ek8gof1KaSirND0WUISBM
qJpPSzOInb9bbxPli7UIVrxVdhinMcMPeHx3wRIGXYEovujEM0+voi8PVV5fiHjl
R+4Ldgb02i83wIGqa8NDgOVpcPpp+R75Q1KVLuqHgIRfmlsiEwWd5jlxPewguIdR
VSeJXVK3CMCnsPP5E1xzgcjJ2OqQB+Zu+Mm9m5rziKtf+0eYRNTtYX3dzqYa5jIL
lvBIjnU1rVQ/7Sbma5KVfEE8ic6/LGGD7cGQ0fcvJXvP1O8X+JOq6+gwOQKw/p3j
xth/sXAdCoWFKWrVwruACRBmi9HuGWYh+hFzxFTVAT+psONPa090Tci7/GHRfrwt
N+S0BX/r17pRuCFecvcnGvPNKiKYVTin45979qrw0fCrRoGT+ugQWIyeXGMWEufh
qyDHV4vjWyElGw5zmU4txGBHp8yfk53EoyMhG6GUiv87VzTUtfIu7kpGZMdi8qvQ
zqBlk6V/YTMxedZrExzpz746plDMKdXGzNVCYV76AAeOYZSEN1Mz6U2NSioSUYu+
e0jeMAe5M5uN4Szp4fzKSbacFPxcwGPw9AGPw5VXqCn4fjCTTV1JZknwxul+UMsf
z3/G8oZe+tQBntOBLpe7zUMSd1qLhhfBPMC8+HR2h0tHf24EEWqKNr119xixExLz
hJccNB3VtsIW6eWYUbS+T25d1VGN4Nm+ju8L9kHLoMkY3OcSORS30d/OVOAc7clq
h0c43TDltqBkjI8mM8dsHlf/24NX98UC491cEifxmQnxgIdJEGk32/6zQvnKF1wl
AKrcYIKNz8Ebglo3h21H4mjRkdbg8BHKHwuDeBsTYAVnYqfDbk5XFST60p4FCM/x
9VjTfJYskI8ETcC4uB6D6Jbu+FBUh3/EWJrQ1N9Fm/WaBJUIIvOaY7ieZrSNgwme
0fJs26nYqxNZgqnIxWkBwFs+R/fULzPtcImmp7SqhHpMSt28gIj0zGFDxoG3zRKy
qoT2t0AmTf2IQXgcYztL5o/wymSUnvjdasQaXB6lAmSyUwDdyN3+TV7Q+2O0rKi+
C1yFghcXYi2KL4/uMYIzKCE4tMzNSTqEVPRPsDlODJQQQ3USsgb4Jjcle85NuZXK
1WKEHgIHPtk3+s21bor0zIvDNpJOlIUz063IMIVyjJAS6E/S76HlT2WPR/tIOnvj
UsNVToaYELKV9evZHX4Jzev4QxWgw4EsANkNYrwXfYOCo4M6uH8gvuN5gEAQlhvj
IpZ9NA82SHjyTAA/5spDh4CUMFHrN5g2E2nRCwV16+lcffWzc1b7OE3J2/mgCK8l
mttc3dcGtoKYEQ38oVaZksaT63oejpQ+jiUhMS8QMGQGQ/mzJk8s3OcrR6ydfhb/
jf/9N4MEVNyMlLcthVCOKi8+1BzSVvjyCwgSMlLnxbgKK4D9MFwrD6cHOevbBlDD
4hIGpjnrxI57ppY2TgaAIArqH2iacpWKQzJFduNn+1FhDL1UszCifSg3ojEX+P+Q
IqPh0siQ8vUe9oETola7cvoBFY5YC9/1n/89uEl8V5lxjOPmKTTd60fHgUMHophA
yFe70YRxY6iPhtyycuyOLnq9m/3lenrjdV7hlX+aUaQHial8+wzkjMjBvsKpmsAU
dhZqARduI+ynwYledQiDt5SELWg2ud7cdAO8GLCpEobrODOmRwBykfDzgEVd6ElR
Hxvw/8HRoGtIebmhcvSikTiDEq2RzgT13gMubnMODsQPyRCFllKlq0SdNsiUCSGU
/IUufJHH5RecutiRgXljP1tHbtx+LwSJgmyY5VksqR5C837Ig8jrx353PmbNhWlr
JIi4WWxgVt2R1smAYxzSAAtKQCBkCL32Wsh9pbpZDtCB5oaGVO7zGrK1sFXU9PoT
p8s7NxoUeH1hZcwfo+DScarrVQR5mzsMZ0H8vUXa5r0GZqFTI79wAiZ0MflfnwIa
lB7VQjL3mtFY+EBQgaEQI41M1yWdAuw2L8mf9RUemXZLqY39V+Y5CAz7qohzsQ07
2T/zWqihR5ehtehh7/OoKaVGwA4CW/DK/Xfv6lEaNuJRDnrI71rQF8PFUkKCP3I7
6Tv7p28Dl//k4n78pbaj1d1Vz8QLf2pQLvBxeE1Pi2VoEZQvWAULjKxkejuIkV71
DjlTKSUbG/iE0NMWd1EiYzLMmNjuQFAqqFUvwpY4Fc3XpL/SDrxVZ3F+u5gGEuJC
CWUAPl/EwWBjlzsjgm22fpahkfTtImP7TACac+dm+pdEVFSeTfqiiq8REn3jOR1L
qG0y3BbkFFP/VNKJ61MlfMpjlsLF89a06PbvIYrenq063PstCmNnR4Jl7/dUxJX/
DhdybiCzl1ugz2NcHIiw+KeeTWiDBzGWehMRMBhMsnC3T9/EYGEOcHlT93NVQb8/
iNsnI7rOQqe0q6+JNnS6voRuYlMTS/AKRqtKwP/H/JYK/cDPgAy2PWCZnkKeAnzT
E68r8OqL3ohKaUzKv2fiaZw8EubO4wplb+lXV6vctAfj5naOwPhcTjvCRtEOuOsv
t+Hp2gNNMElc7ObP/Yrl9fRFhXVbcstJvg+iKayGJzIcXQ1/0HedQ+zhc69cCtOz
joBYviN1xnAdTvev8MtTUnlcnKMZNvz1oL5JL+4GNVotQsgXWmipUyfwRcp494aU
Frn9Ximj2O7aGktyFm3z9ZhjYe4WbY174RdEZnuEkzpPa8Qf+mjdojkwLoYRelvr
s8fQ9lPfywI5VJFEZJWgHlK70FtzYAIcjnBvU8bSvhz0d6dD0WLm/vT2oqBgpyjz
tkrGhvbGaxZ7dEaTZzk+ahjWZrw4NiWYKdDirQNIZtMuDkAxi4kfCmY8o97aLSg1
MMlRMr9YEeKM7HoUnh6KOhy42005R/ldYHFFNSvsbzfJUcIpq8lM3TE3+SKXGUi9
z6nYUJc/Gj7JN7tENYrtiMQ/MWtlyy04RjqO7bTbyWiHt+LsZC3ptKBjfqVHUFau
ICDYZOzAwcNgC2TsOslrPGdW+D+MHmaB3yaw6Ncqz9motwUPEbl8XzfiNY+t0rx2
hEjHgLq/MSLpr7H9KELmcIEWYUQLoCSHXOC2haYIJA/C0XaDEk2PvrwQVwhmS+u1
Ai4EECY/TbabK4zqf8MIVdNTfJ6IWrjQzeaWf650gPfWMdZoRUUwNvttpGYwNdjm
UTNnhzOM8/zSogPsMreAqpxsrjdxeB/xGOwbRTP6gxyNrnwybDTgniJiH3VnzEYA
PdUsPwrS0/T74WEuH9KtUtiC6w6LCYxHhVNsXvKoUYr03xeh4lKE6ymO0d6NEGXk
hWfSSrk8wQ890eCLu56rWASoEc+TmTnO4RSI9zvR4MnSvI7pP+rFU15wbRUwyXjX
fwqD+4gJIzzlzs5tHK7zgdS4hDLL7FZL7ZKQgihWogXsvnClz3Y6ASXW8gvsK1Eg
XWGQuwwXrfgLuNSF6QKitsB3J3V3744593znKcbd5S3irRVmD5GkMey5FfOxs3Ig
ouBrLj8wu0ZMjaRWUyInGj7d/XoZwg/opJszY62BKu7dVSbfhs790Tfu3c3VlvWO
QfOAvPxWCUwy9MXefXFm7M3xyYM4PHhl4jSBeLqf+wDuIuHu/VZ9btn71pj7OOCb
DgydudeusXmAsCrlWasQlNUgkF4LCw2FssBwiE7bSnP7NsyO6khqcGHw0Ekm4cS2
BMvrzO//hdqRK5liopZULVe9arp3I/nXMB+7GzAtgKuqKABHWnxldDJeqJtnEMT1
2J61K4PwmNY0WXUI6eTSmv6iE8uxB+Uq5FY4ZNYiyxJBcWjLMTBm11JyyfUd5cnz
yj1XXTDK5fN/d53FlU6pOh/jsqHEbsAYeTSox/N3ZUROV7R5+wvsygGfiKJWVsPA
JqH9OHatePIZiqxGWH1bFCDpSZndklzXr7djclto4UZsw3MTXTVvWCVI63Q6lxg3
QxOVGcmjc7ZQ4Fb7UZuaXKgbbm5irCkyN1b6fYa4jd8ot/jU9/N1OoRePeddfOIQ
xvPDEuipe081imv1HcDe462I/ZU+Dgk3FTkSFF8ZmuQhpKBesvvZ0b5jX0hZi4+j
xTcq2rMFM00QvXBVwhUjf6Qg80O7gU1PSCywkHBQDlJskKGnNXQbS5HBzuFjMK1O
6nFw+P440fxqtdJipSXJBvzqGQsxB2s65ZGDdpHH29Jgw5MGWcxKGQf+3DKK75Lq
ZNVDFfvXXSw3QN9JYzUSMVx03qn2LJgcNTLa9GPSncGZL1PbN6wxgDZwbWpOQCpg
a3QHvUUME47PTXEyYCCyXNHgF+hTwawY8lLaMdloYoHmYnhki3UYfj6Kb/dQl/ZD
492gontUEkf9ZhUR8dzKTjH2thaglhhuiYyZDzBn1eBDn+LrR2ECQhs0DlcgZAhK
7XEVH3pDAOgAzn9Xqk+iAZAXPbwS5qR5/5yLd+QANh4wOvPNfq8z8+kiFDgvhx89
`protect end_protected

