`protect begin_protected
`protect version = 1
`protect encrypt_agent = "Anlogic"
`protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-002"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
XIeluV+BBYty+J7SK9a3UGm2jxmeSdR0RtDrPQwHYwTFmsV2WLyVjLeRrBjqwWNA
Slsikgt9UFdU6SADK5ryV3evLC7CzlUI9JwWhDv0XS7FC8XQdcL/yarXrxCeHh5D
iIckTpT2Jz/ogIAr2H4gCcERorIyyNu2zPXnbNHy4uc=
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`protect key_block
op0+bpgNdc3mCRGHraeBH9WzAIBR6TYlhZe1Rus4zad2Nf23vKw8nVKFYgJKNlJt
+ZrtWqK8dKEJHMhv6WNHi5DsfGRC/tdjOXfaGZFTMGebB1FgtRSSjOEi0AHpjINU
Ljwoys2cddd5tATi31wz/OIAvHvoipBXTXSV1y8zaXjh0OHH4wxicJORYRcJW5Iz
ZtOmX6zCQaMLNDs2NvePYW4IbyxhZVpRFawjIm+FkLWasSV3K7k7dTwKUNtDEYPy
atEbHcM1iELBClMtTYZCzYIxrlcbrqPr4VQhtSh0szleWyMMgzjC48iQRlEFEkQn
EgCJuiryP5InKIJ1xr9KkA==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
EBunLZCnrnynvTewsInXGtwiwkUwfPzIH/T94xt/KHQi3fRlf7Fu9WGCmXcoUYrC
zf74VrXiBG8ArK2gHt4d81meNaZ+E7fsFbQgbhKUFGk54VXZvCUGjRywirKf9C7E
g4pCuHWen5/RUyx9ZTsMT6Z5DdmMLrvzKSzc1wAaMXQ=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`protect key_block
m+I2UcvClJYsQMLIi0KDODyyYMTBqbOwR7iAduXdKcIUFivjo7KGp+M0a8vrgbxd
3GgsK7epQqORzX1XoXnIeeuBVD13mzKW4INDzXO28XYlggBq8tzHSBc662P84R5R
S82GThwfMbffQjRbpSQnqa6GR3Jz+yk0iSiROU/DjnT8H9xtDbvwf51F1quiU7xX
aQp35gbb417P49x3AYyfC9aEl4LuspkxDE/4WiBBF+YBZOBFEqOF1rNXf2YP6+Je
ko0Qm/qRVz1gRxqpQWQPoPrimKZjxN/1s+QjD3fk83m0lS8ZLc9Tn0Zpz1SyP+Nv
d3HG+sZQLE3t/TwPYbb06Q==
`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
AmIwFgczimbwCaNWVM8TeOmJqQxcG/YJncBCTL2Um0QqtjpDoXVkuDL0CYsfJbez
NDnAsqjhqi6AzqnaE4myE3dvyzN+VbaFDZ2MJFpo9l01q0vFkDZZED3Lvhx+pllI
1fnYedLur6Iy0kb4hgHaewy7twBpWlvTWv2VOOe/SpA=
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 4000)
`protect data_block
S01Ib1g4Zkx6emtZSHJuWC0wUGm6aIOdHrg5gJPwP/EKryNF4rfgj+9pw2cJY5nN
lpwxB+oGdwJd+4jYdMhTC6bJIgXpq24c5H68cnnJTfduTKbD2zcjh/Wd0AUnL4+c
u99foCh4eihfJtgkF4IWD6MKu0C9wdVLdg1IqyJt73LZQKdVE0VkXYuZJH6VYvjW
a+uneaT7X9D/yW+vZcy0z8vEA+eZ180163MVJrz/X0eQKM3QlbjM+s5+ECaF9Zix
3vstNFEoLTzuXHo/C6uOrQqmwqyI63TREoXsowVWkQJCqbVzELleV8TZ8qYiGCHU
CD5GnXK4mfCPwP6OWvgMdw0CgDBDwG/GAlMgTByVbrFNQmdc4Kv0ARLgpCVsvIFx
MyowejCeTqcEMUbDs4bhn2iodMF37XVVgJdw+1oZV/PiC7/mXM+zwAkqzisQw2Ve
vjJ516gp/Xyt9XDjLYu4nEzkXYxSduu7VS4NqFMbYSOKV65lHdK3zxwMg/V3HKE0
HMnkchEfsQMQeva9xvGbmrJOUALFInsM2NPlOGmP8V450SOazb2yFsKky2sptfRc
VKQ9r+BpsWUD8C6y2WG2/C22pNs2Gb4Lbw8O2MTDEOzWl7wCoPYQVhbcBdP17ilF
tBhQziLRtUnWJntutwTHKv9UVDrpUiXTue+8cls09WzH2V+CLSeup+p8K72baTgs
l8PDYY9mGypZo4p6nqTgA1tSo2WkSUe/UexKH0S5u4jRe3VpPxpuoeVdZ9lWKbFJ
rNfxqP00VWaIbPgnZLp2XnvfxWirBumI5lBeeZix9dAGTmZnvyiqNUF/CtbVatQP
6gnoDecZEnAtZtT2jO1VoWyZKbiyUVXS1eNzsHBcB7qlJqPmElZ45phLjzdZ2DwH
lYfuON8RJm6sSqcEE5TNc34+qSzO3ggCZR4L7SpuJifkCA0xMSrgm7PEEh1rCJKk
JjJWvTIGT/Eijs5ZqLT5w0T8U6mdhw8CwBq5BQamgIpkCxeHpsAb7oL7u7qMVCG2
4I/FqkONOf06IUie7UIYuyRDNh7zKn4jmlC7WwNixrIqWfss96dm1zLhbMuYTyZ7
ULjEi1RmgaGqGNJsvOJeFrs7DHdEy+77jBW0zrnXFPbfKVJ5+lOqB74tvFGgkTf3
4qpfvZ/l+rRdRSlVsWpXhO/tIRDYpVSGZcH/17PKBNI/uuJFfWjjf4Jas1aOZKnG
piTiTKGij+lLIvalkxOI0RyX8aD1exXBnhFmUlFBMLSulMLJoi24OMqoROFy5ozc
FY8ZgFXbFv8o5dYekm8x9Uxpoq4Yfqy9z67Oo8BhLD7/yfA6tsM1LDJDzNkIAQaQ
7hlVGdiehcv3H5A5tQ2dP09srrL3Uin1i0v1aOz2E1qL0qrOLnH6wbygY7B4M1V8
VmFZS+l3ZFD/gQzLv0PnPkz0T5H3pMSTiLMfd+dNlCQxJH6R8a+tEx9+0F4AKPie
sdfpzfFjpYaFklF5ItBrlHB9LLCQWHSIw4bIED9NjJ6tC3ACxKeij2eEneWf3qem
XJBnP0IsKmiIhij23L4UXsTcd+SoOIvtZ5TNKsjo7p2/zhZylrObeRDvD1UTqoQC
GplA0P6woOZ2oUw9aL8GFKXmSoIt7ZTZ3TIp4ZcUq51kdhPUBoD7SYtzUYaUACG3
H5Mu9Hg1PXwP+1yn4GIEk/KYV2Md3e9WLNPbtyE2pDImNWWkhKu3Et2KEmU6H6xd
a1U+2wLmdB/VKdPDWMb8LQLaKF8ovviYLFN1zIRuD5hyrrgvtt5aLPGMMAGmLvDe
xefvormLnW4HMtr+yylWpf2FnlQiIPbr2CqElzqH8xy5arAI5SzZ/n72wV8ivFg7
Ym2yz22WuhAfo+tUipzytERPoJKswM1gXAGHNAPIrWVitoKV8I0Lc+Et3vkcczBk
2kPPAPllDKxZmGUKbFHX0QII0UpNGt+Woc5dVTA1fhB4aaLUnAz4kZZpaMU26PEA
Rylepfp5BwHhkUAg4PQx8EtM+n01r84sH6FYsSEpVJ/aTHelcxUpooP2KO6CIPZK
YQlIf9FzbaXN+9eBLc7Wt2ITR4nzurQGT2xUPySJB9AnAQErRgcPjOHXjKLoQsOB
RDDztCvIH0gXoEFiq0rCY0Ehu7KRin6jcux0s9TmoNmDd8fB7rtYnT6IJvbr20DH
jb3gJLUOsaQp+kAQOWubYjv/pcFeNkc3I9czu/0XFRt3lKYcM6sCxvBflP6fTpVP
m+JWXSmwZHPhfxVngZDFA6VOMAbJ8pi0XYjIyqlftEr41acIBs3CjvN6Ll7rePyj
aFa3raV+qAIUx32n1CF+y6WjSGx+T/nerkYBU2ibCFaTIA4bWEOalboU4gR3aONA
rtY4ohJoQsYVh6Uaw9IOi3R7m5s+hQb0Gc6D99iU5ljAotNp2/GhT7qeGNUMmea7
lzsG9BddN7aMiMFdQ6qPRet6qi2dO4wfs4zQzPgh7CLHaZz0Sk51u9fJiGf4QWJG
Zcf19Fu7Uq23CS9DZSc1tmx//z+W2lc5dw4v/LDCPonLavvHgSwaLfm/jp+JbuRG
w1WA0n64jsbs3Kib4lShyOrw5U14mRjT+HH2RwWGA8eMH423evfI9rdXGK0//5Wx
3HRCmnIt4QKw0vrjvOtDhyRcFT7oTBbaZpi0fIDIr1rY2Uja7mljTwhbQd8ZjLo9
HXwzhLDyTUaZqi5mtLkgsIMLmghBBrhuH9penDY2sfkLd60TNR8M6cejafZaASAp
+OJOZHknit4j/62JC8H3xRav2yU+Mk3NPUUO2YzUSB4pPpp40kQjnqbQeEo8QQIj
ulK+MYzDkdIEAQteXyr6ZLYKKXIARPYlftG7Q+SmI6FFWybxfhQmrIMUzdjo8wWP
WB3Y7qqHBlLUag2fSHg2nZ/rXsTKzaeKlm/PzkE5pItqVubc70p8ylXkLbEzqXLg
T0t8w660C05LUh7dj4vhuL4tJIMkEkV94JERP6EjixOzouiYMRA7ux/OLZpsFTa0
9WnBzv6n/7sJIwgFstHgkF66o4Z7HJPYFvyD9QVxS4YNp6cW2Pssz/Bak0gSTUHt
gDBZEbgPjyhxvebz+OevG6Z4CYBxDEXM2452GrJ3sQn1e5vHG3mgW0CEw9tN33vz
gn1oRQYKO/RemklGMShfLgI2A98xS7FVOEHnl4D+bBIxxe8y/7I2LDRdOBrlmCsu
okkAAmZflOh9Yi8ASSLo5waYj6Izdu7m7hMeWzsC6qV5zlLTofBwpdnKRSyIPGEJ
6nk880FdjjYSPx3v+bkQKMkivUFCD86z3cyBD3vXUPvcnHSzHzc1Yliy73KcDlyx
K3Ilt8XDWAThIRIhBfstqkqhM37VMMy30xIXfwjbhDDDgHhpczpyZuBddFurDznF
n5arHRBYLRgVw9JU/1H2jJTy0lFX22I1Apv8hcrPkGI6AXkOF/T33Vsu1WklR5rK
FRFZoG19ehpN2el7Ldf17o3Bm/8P+8m6wxYMNVEHWYY9VHsZRxAzwXUCu/Q6X9nP
cKFfO4Sn74hVfRJXQaqG01VIFWtTdUKjb4scJSA/ntKNrZpyRuys80teX1k/iYKZ
oyUonoSOuHTsErTMH2mvdR3Ti7kjQocRwqYm6prMfRRZ21z7zs8L4XyaNlrhZ0t/
Q6NQnPzbIa1UR/8yNn7wSFfCEMAA7J7PTjEhidkRGF1mHtrWCMHmpRi4ExRRuRUM
h+DPRuOqB6iopNtjVlJ1gaj704QSgFrbgVgjs+gUi4Gqf3RUGvxGz9UymGCBS9+a
lif7k0omRa5BrpYPdciq+myKzRxOy2wdMFh3nCCOznFhOjo4ZfGkGaiS1Fv37oXy
aL1Q+pLr9K6xwBD4sRgrXWz/s3SICs4jts5b24jrqMXZkeSTpMINTV4NhkwpM1GA
p5rGDB5oJXpunAxDVJvrpqfNqURr/VXHB24tbkHa/91yj6kX2FS8koBURPlM+LiV
SslNHa7vSw0QDJqgRQoRUpGzseJikK7PjvdH/j4lvCyif5Q6ymkhfHrAw0AJIYsk
yBCx7PmRDHtahvrVBW5h5erz84d2+5AXRM0dsghl4sFONrXXHVMD4tEtDqsO/9/3
IlEAIWdnWi7uldeVP22pcR3Y5ASgYJjew4LhTwusyHuPllSrpRmLVEv3rF6MY7//
tqwQToRlgykM0pHawVwDsstwESNxN71reNKnQDDM0/EwV+wUBZ1fWtZQAr1ZeBPx
EtLFD7Jcci9azGAIcD6ApxLy2NFxuw3hdf3Kyy4ZtsF6OKQG2Jm5EsnU3O2KYGt6
FlsHyI4rZ8VxYYnzawDpxUGoEje3+OTiLW1zPrXUVZFp05RiPjILKtuB567vHxEJ
4djdqRlQBwJFXCqbbvy23FN9X/jXyhhwK39MyYtEKW5bxjZS98/txnSFSPbn4Jw+
f3pLZ6UMnq2ci4TDWfo9EkMa8xJLL9LL1kZEglF2Ro8eYWQkcHTU3e1nbmmpMf1X
jNeUcNXVftd7f11EbjdIvScH+Z8pvyVboMysgXp9mU+uj/8T1r1/BAvu08NpRabT
+TkjvN7eDVuJ8vGXVdD6sAypH87Yl+5rfOYFgK4TkX6y3xKDyTR0DrU1Ai06ZzIl
QZpnsYC2n7id6Ge3T5BJKaLjaOxH7RwfSnwh/3ozgCtczAeIk6Te4pRUda4I7ogC
LZhUbpMyLF89v6/ZozfhQrxpN0bh8Yz0NKESt27Vtv1Do3mlFWWYx5tdXRTXn4pZ
N6xBA3+K2tejLafqLvR4elTQS4BYpkGKjwoxJW6fMJ0AGr2Kz+KcX/6ln7DzhwPS
sG4Yr1RBopR+nDKGwMMUyB8J3F6+zjdeSUJBDMJtljlwH+NIRkggy4GzIyfLNdJI
UNc6uO66sNnK6JVLllpfvlg6TUGn215v8jL+G8oAVsrGF6wUqsWQf+E8TD6Rk5in
NjtleUejx/WWKTyMW9vTdrVdBdjWLpvjukmU51ej/xoA/9YkoRjBWG5SSOyoxiUr
oPNyyAj1R0Cbs/rUZ6kZzDLM5T7L2G538hOZjANxv78KJ+/CaOizUWLxopNoSXyu
z6usFV3nO8ZxLYWkZI6thZ8IkuhM6GH5JFCTc+1dKfeViETlPaYY3giq869c6cq3
UHa/L9rMhwMhQjHWNxykh6K1AqOx9TKsWXWx5dX633fiKisReZsdrICp5Q4s5eNN
SvFVEjzrraK957YJdTq9jgnwtulJ50bzNuvIYn8PMSfKElCqqZOtbYZ4pyVOc8Z5
gO602RdUieNG/8smKN32cl2wTOAGGen4UyFg/o7OsIjRUSd7JPSh3vs1uZRsKUqL
PF1adaJdJA1Ur1lDnITLjw==
`protect end_protected
